module main

fn main() {
	cli_setup(compressor)
}
